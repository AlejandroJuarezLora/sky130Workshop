magic
tech sky130A
magscale 1 2
timestamp 1718324108
<< error_p >>
rect -29 127 29 133
rect -29 93 -17 127
rect -29 87 29 93
<< pwell >>
rect -211 -265 211 265
<< nmos >>
rect -15 -117 15 55
<< ndiff >>
rect -73 43 -15 55
rect -73 -105 -61 43
rect -27 -105 -15 43
rect -73 -117 -15 -105
rect 15 43 73 55
rect 15 -105 27 43
rect 61 -105 73 43
rect 15 -117 73 -105
<< ndiffc >>
rect -61 -105 -27 43
rect 27 -105 61 43
<< psubdiff >>
rect -175 195 175 229
rect -175 -195 -141 195
rect 141 -195 175 195
rect -175 -229 -79 -195
rect 79 -229 175 -195
<< psubdiffcont >>
rect -79 -229 79 -195
<< poly >>
rect -33 127 33 143
rect -33 93 -17 127
rect 17 93 33 127
rect -33 77 33 93
rect -15 55 15 77
rect -15 -143 15 -117
<< polycont >>
rect -17 93 17 127
<< locali >>
rect -33 93 -17 127
rect 17 93 33 127
rect -61 43 -27 59
rect -61 -121 -27 -105
rect 27 43 61 59
rect 27 -121 61 -105
rect -95 -229 -79 -195
rect 79 -229 95 -195
<< viali >>
rect -17 93 17 127
rect -61 -105 -27 43
rect 27 -90 61 28
<< metal1 >>
rect -29 127 29 133
rect -29 93 -17 127
rect 17 93 29 127
rect -29 87 29 93
rect -67 43 -21 55
rect -67 -105 -61 43
rect -27 -105 -21 43
rect 21 28 67 40
rect 21 -90 27 28
rect 61 -90 67 28
rect 21 -102 67 -90
rect -67 -117 -21 -105
<< labels >>
flabel metal1 s -45 -28 -45 -28 0 FreeSans 480 0 0 0 D
port 0 nsew
flabel metal1 s 45 -29 45 -29 0 FreeSans 480 0 0 0 S
port 1 nsew
flabel metal1 s 2 110 2 110 0 FreeSans 480 0 0 0 G
port 2 nsew
flabel locali s 0 -213 0 -213 0 FreeSans 480 0 0 0 B
port 3 nsew
<< properties >>
string FIXED_BBOX -158 -212 158 212
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.86 l 0.150 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 0 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 80 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
