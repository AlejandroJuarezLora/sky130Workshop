magic
tech sky130A
magscale 1 2
timestamp 1718753713
<< error_p >>
rect -29 90 29 96
rect -29 56 -17 90
rect -29 50 29 56
<< pwell >>
rect -211 -228 211 228
<< nmos >>
rect -15 -80 15 18
<< ndiff >>
rect -73 6 -15 18
rect -73 -68 -61 6
rect -27 -68 -15 6
rect -73 -80 -15 -68
rect 15 6 73 18
rect 15 -68 27 6
rect 61 -68 73 6
rect 15 -80 73 -68
<< ndiffc >>
rect -61 -68 -27 6
rect 27 -68 61 6
<< psubdiff >>
rect -175 158 175 192
rect -175 -158 -141 158
rect 141 -158 175 158
rect -175 -192 -79 -158
rect 79 -192 175 -158
<< psubdiffcont >>
rect -79 -192 79 -158
<< poly >>
rect -33 90 33 106
rect -33 56 -17 90
rect 17 56 33 90
rect -33 40 33 56
rect -15 18 15 40
rect -15 -106 15 -80
<< polycont >>
rect -17 56 17 90
<< locali >>
rect -175 158 175 192
rect -175 -158 -141 158
rect -33 56 -17 90
rect 17 56 33 90
rect -61 6 -27 22
rect -61 -84 -27 -68
rect 27 6 61 22
rect 27 -84 61 -68
rect 141 -158 175 158
rect -175 -192 -79 -158
rect 79 -192 175 -158
<< viali >>
rect -17 56 17 90
rect -61 -68 -27 6
rect 27 -61 61 -1
<< metal1 >>
rect -29 90 29 96
rect -29 56 -17 90
rect 17 56 29 90
rect -29 50 29 56
rect -67 6 -21 18
rect -67 -68 -61 6
rect -27 -68 -21 6
rect -67 -80 -21 -68
rect 21 -1 67 11
rect 21 -61 27 -1
rect 61 -61 67 -1
rect 21 -73 67 -61
<< labels >>
flabel metal1 s -44 -32 -44 -32 0 FreeSans 320 0 0 0 D
port 0 nsew
flabel metal1 s 44 -30 44 -30 0 FreeSans 320 0 0 0 S
port 1 nsew
flabel metal1 s 0 72 0 72 0 FreeSans 320 0 0 0 G
port 2 nsew
flabel locali s 0 -176 0 -176 0 FreeSans 320 0 0 0 B
port 3 nsew
<< properties >>
string FIXED_BBOX -158 -175 158 175
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.49 l 0.150 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 0 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 80 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
