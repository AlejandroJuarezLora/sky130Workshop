magic
tech sky130A
magscale 1 2
timestamp 1718320476
<< error_p >>
rect -29 308 29 314
rect -29 274 -17 308
rect -29 268 29 274
rect -29 -274 29 -268
rect -29 -308 -17 -274
rect -29 -314 29 -308
<< nwell >>
rect -211 -446 211 446
<< pmos >>
rect -15 -227 15 227
<< pdiff >>
rect -73 215 -15 227
rect -73 -215 -61 215
rect -27 -215 -15 215
rect -73 -227 -15 -215
rect 15 215 73 227
rect 15 -215 27 215
rect 61 -215 73 215
rect 15 -227 73 -215
<< pdiffc >>
rect -61 -215 -27 215
rect 27 -215 61 215
<< nsubdiff >>
rect -175 376 -79 410
rect 79 376 175 410
rect -175 314 -141 376
rect 141 314 175 376
rect -175 -376 -141 -314
rect 141 -376 175 -314
rect -175 -410 -79 -376
rect 79 -410 175 -376
<< nsubdiffcont >>
rect -79 376 79 410
rect -175 -314 -141 314
rect 141 -314 175 314
rect -79 -410 79 -376
<< poly >>
rect -33 308 33 324
rect -33 274 -17 308
rect 17 274 33 308
rect -33 258 33 274
rect -15 227 15 258
rect -15 -258 15 -227
rect -33 -274 33 -258
rect -33 -308 -17 -274
rect 17 -308 33 -274
rect -33 -324 33 -308
<< polycont >>
rect -17 274 17 308
rect -17 -308 17 -274
<< locali >>
rect -175 376 -79 410
rect 79 376 175 410
rect -175 314 -141 376
rect 141 314 175 376
rect -33 274 -17 308
rect 17 274 33 308
rect -61 215 -27 231
rect -61 -231 -27 -215
rect 27 215 61 231
rect 27 -231 61 -215
rect -33 -308 -17 -274
rect 17 -308 33 -274
rect -175 -376 -141 -314
rect 141 -376 175 -314
rect -175 -410 -79 -376
rect 79 -410 175 -376
<< viali >>
rect -17 274 17 308
rect -61 -215 -27 215
rect 27 -215 61 215
rect -17 -308 17 -274
<< metal1 >>
rect -29 308 29 314
rect -29 274 -17 308
rect 17 274 29 308
rect -29 268 29 274
rect -67 215 -21 227
rect -67 -215 -61 215
rect -27 -215 -21 215
rect -67 -227 -21 -215
rect 21 215 67 227
rect 21 -215 27 215
rect 61 -215 67 215
rect 21 -227 67 -215
rect -29 -274 29 -268
rect -29 -308 -17 -274
rect 17 -308 29 -274
rect -29 -314 29 -308
<< properties >>
string FIXED_BBOX -158 -393 158 393
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2.27 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
