* NGSPICE file created from opamp_plano.ext - technology: sky130A

.subckt opamp_plano vdd gnd vout2 vout1 vb2 vb1 vin1 vin2
X0 vdd.t33 Y.t2 vout1.t3 vdd.t32 sky130_fd_pr__pfet_01v8 ad=0.93885 pd=6.02 as=0.93885 ps=6.02 w=5.69 l=0.15
X1 gnd.t11 sky130_fd_pr__nfet_01v8_DAKYLM_1.D sky130_fd_pr__nfet_01v8_DAKYLM_1.D gnd.t10 sky130_fd_pr__nfet_01v8 ad=0.957 pd=6.13 as=1.798 ps=12.22 w=5.8 l=0.15
X2 gnd.t3 sky130_fd_pr__nfet_01v8_DAKYLM_1.D sky130_fd_pr__nfet_01v8_5Y6VJK_0.D gnd.t2 sky130_fd_pr__nfet_01v8 ad=0.1421 pd=1.56 as=0.1421 ps=1.56 w=0.49 l=0.15
X3 vout1.t0 Y.t3 vdd.t31 vdd.t30 sky130_fd_pr__pfet_01v8 ad=0.93885 pd=6.02 as=0.93885 ps=6.02 w=5.69 l=0.15
X4 vdd.t7 X.t2 vout2.t9 vdd.t6 sky130_fd_pr__pfet_01v8 ad=0.93885 pd=6.02 as=0.93885 ps=6.02 w=5.69 l=0.15
X5 vdd.t40 X.t3 vout2.t8 vdd.t39 sky130_fd_pr__pfet_01v8 ad=0.93885 pd=6.02 as=1.7639 ps=12 w=5.69 l=0.15
X6 vout1.t5 Y.t4 vdd.t29 vdd.t28 sky130_fd_pr__pfet_01v8 ad=0.93885 pd=6.02 as=0.93885 ps=6.02 w=5.69 l=0.15
X7 sky130_fd_pr__nfet_01v8_DAKYLM_1.D sky130_fd_pr__nfet_01v8_DAKYLM_1.D gnd.t9 gnd.t8 sky130_fd_pr__nfet_01v8 ad=0.957 pd=6.13 as=0.957 ps=6.13 w=5.8 l=0.15
X8 sky130_fd_pr__nfet_01v8_5Y6VJK_0.D vin1.t0 Y.t1 gnd.t12 sky130_fd_pr__nfet_01v8 ad=0.2494 pd=2.3 as=0.2494 ps=2.3 w=0.86 l=0.15
X9 X.t1 vin2.t0 sky130_fd_pr__nfet_01v8_5Y6VJK_0.D gnd.t12 sky130_fd_pr__nfet_01v8 ad=0.2494 pd=2.3 as=0.2494 ps=2.3 w=0.86 l=0.15
X10 vdd.t27 Y.t5 vout1.t1 vdd.t26 sky130_fd_pr__pfet_01v8 ad=0.93885 pd=6.02 as=0.93885 ps=6.02 w=5.69 l=0.15
X11 vout1.t9 Y.t6 vdd.t25 vdd.t24 sky130_fd_pr__pfet_01v8 ad=1.7639 pd=12 as=0.93885 ps=6.02 w=5.69 l=0.15
X12 Y.t0 vb1.t0 vdd.t35 vdd.t34 sky130_fd_pr__pfet_01v8 ad=0.6583 pd=5.12 as=0.6583 ps=5.12 w=2.27 l=0.15
X13 vout1.t7 Y.t7 vdd.t23 vdd.t22 sky130_fd_pr__pfet_01v8 ad=0.93885 pd=6.02 as=0.93885 ps=6.02 w=5.69 l=0.15
X14 gnd.t7 sky130_fd_pr__nfet_01v8_DAKYLM_1.D sky130_fd_pr__nfet_01v8_DAKYLM_1.D gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.798 pd=12.22 as=0.957 ps=6.13 w=5.8 l=0.15
X15 vout2.t7 X.t4 vdd.t44 vdd.t43 sky130_fd_pr__pfet_01v8 ad=1.7639 pd=12 as=0.93885 ps=6.02 w=5.69 l=0.15
X16 vdd.t36 sky130_fd_pr__nfet_01v8_DAKYLM_1.D sky130_fd_pr__res_generic_po w=0.33 l=1.65
X17 vdd.t21 Y.t8 vout1.t2 vdd.t20 sky130_fd_pr__pfet_01v8 ad=0.93885 pd=6.02 as=0.93885 ps=6.02 w=5.69 l=0.15
X18 vdd.t13 X.t5 vout2.t6 vdd.t12 sky130_fd_pr__pfet_01v8 ad=0.93885 pd=6.02 as=0.93885 ps=6.02 w=5.69 l=0.15
X19 vout1.t8 Y.t9 vdd.t19 vdd.t18 sky130_fd_pr__pfet_01v8 ad=0.93885 pd=6.02 as=0.93885 ps=6.02 w=5.69 l=0.15
X20 vout2.t5 X.t6 vdd.t9 vdd.t8 sky130_fd_pr__pfet_01v8 ad=0.93885 pd=6.02 as=0.93885 ps=6.02 w=5.69 l=0.15
X21 vdd.t17 Y.t10 vout1.t4 vdd.t16 sky130_fd_pr__pfet_01v8 ad=0.93885 pd=6.02 as=0.93885 ps=6.02 w=5.69 l=0.15
X22 vdd.t11 vb1.t1 X.t0 vdd.t10 sky130_fd_pr__pfet_01v8 ad=0.6583 pd=5.12 as=0.6583 ps=5.12 w=2.27 l=0.15
X23 vdd.t5 X.t7 vout2.t4 vdd.t4 sky130_fd_pr__pfet_01v8 ad=0.93885 pd=6.02 as=0.93885 ps=6.02 w=5.69 l=0.15
X24 vout2.t3 X.t8 vdd.t38 vdd.t37 sky130_fd_pr__pfet_01v8 ad=0.93885 pd=6.02 as=0.93885 ps=6.02 w=5.69 l=0.15
X25 gnd.t5 sky130_fd_pr__nfet_01v8_DAKYLM_1.D sky130_fd_pr__nfet_01v8_DAKYLM_1.D gnd.t4 sky130_fd_pr__nfet_01v8 ad=0.957 pd=6.13 as=0.957 ps=6.13 w=5.8 l=0.15
X26 gnd.t14 vb2.t0 vout1.t10 gnd.t13 sky130_fd_pr__nfet_01v8 ad=0.3886 pd=3.26 as=0.3886 ps=3.26 w=1.34 l=0.15
X27 vdd.t3 X.t9 vout2.t2 vdd.t2 sky130_fd_pr__pfet_01v8 ad=0.93885 pd=6.02 as=0.93885 ps=6.02 w=5.69 l=0.15
X28 vout2.t10 vb2.t1 gnd.t16 gnd.t15 sky130_fd_pr__nfet_01v8 ad=0.3886 pd=3.26 as=0.3886 ps=3.26 w=1.34 l=0.15
X29 vout2.t1 X.t10 vdd.t42 vdd.t41 sky130_fd_pr__pfet_01v8 ad=0.93885 pd=6.02 as=0.93885 ps=6.02 w=5.69 l=0.15
X30 vdd.t15 Y.t11 vout1.t6 vdd.t14 sky130_fd_pr__pfet_01v8 ad=0.93885 pd=6.02 as=1.7639 ps=12 w=5.69 l=0.15
X31 sky130_fd_pr__nfet_01v8_DAKYLM_1.D sky130_fd_pr__nfet_01v8_DAKYLM_1.D gnd.t1 gnd.t0 sky130_fd_pr__nfet_01v8 ad=0.957 pd=6.13 as=0.957 ps=6.13 w=5.8 l=0.15
X32 vout2.t0 X.t11 vdd.t1 vdd.t0 sky130_fd_pr__pfet_01v8 ad=0.93885 pd=6.02 as=0.93885 ps=6.02 w=5.69 l=0.15
R0 Y.n0 Y.t8 1150.05
R1 Y.n8 Y.t6 1149.41
R2 Y.n7 Y.t4 1149.4
R3 Y.n6 Y.t9 1149.4
R4 Y.n5 Y.t3 1149.4
R5 Y.n4 Y.t7 1149.4
R6 Y.n3 Y.t11 1149.4
R7 Y.n2 Y.t10 1149.4
R8 Y.n1 Y.t5 1149.4
R9 Y.n0 Y.t2 1149.4
R10 Y Y.t1 117.392
R11 Y.n10 Y.t0 111.635
R12 Y.n4 Y.n3 6.02208
R13 Y Y.n8 4.35576
R14 Y.n9 Y 1.48734
R15 Y.n9 Y 0.833298
R16 Y.n1 Y.n0 0.650756
R17 Y.n2 Y.n1 0.650756
R18 Y.n3 Y.n2 0.650756
R19 Y.n5 Y.n4 0.650756
R20 Y.n7 Y.n6 0.650756
R21 Y.n8 Y.n7 0.642604
R22 Y.n10 Y.n9 0.476616
R23 Y Y.n5 0.340334
R24 Y.n6 Y 0.310922
R25 Y Y.n10 0.00593478
R26 vout1 vout1.t10 62.3383
R27 vout1.n6 vout1.t6 44.8719
R28 vout1.n2 vout1.t9 42.8569
R29 vout1.n6 vout1.n5 38.6225
R30 vout1.n8 vout1.n7 38.6225
R31 vout1.n4 vout1.n0 38.6225
R32 vout1.n3 vout1.n1 38.6225
R33 vout1.n5 vout1.t4 5.71315
R34 vout1.n5 vout1.t7 5.71315
R35 vout1.n7 vout1.t1 5.71315
R36 vout1.n7 vout1.t0 5.71315
R37 vout1.n0 vout1.t3 5.71315
R38 vout1.n0 vout1.t8 5.71315
R39 vout1.n1 vout1.t2 5.71315
R40 vout1.n1 vout1.t5 5.71315
R41 vout1.n2 vout1 2.42124
R42 vout1.n3 vout1.n2 2.01553
R43 vout1.n8 vout1.n6 0.537265
R44 vout1.n4 vout1.n3 0.537265
R45 vout1 vout1.n8 0.276235
R46 vout1 vout1.n4 0.261529
R47 vdd.n26 vdd.t34 909.881
R48 vdd.n12 vdd.t10 909.881
R49 vdd vdd.t36 613.304
R50 vdd.n25 vdd.n24 525.279
R51 vdd vdd.n1 324.118
R52 vdd.t10 vdd.t39 210.643
R53 vdd vdd.n10 158.381
R54 vdd.n25 vdd.n13 113.942
R55 vdd.n1 vdd.n0 112.733
R56 vdd.n13 vdd.t35 110.085
R57 vdd.n0 vdd.t11 110.085
R58 vdd.n24 vdd 74.1861
R59 vdd.t20 vdd.t24 57.8685
R60 vdd.t28 vdd.t20 57.8685
R61 vdd.t32 vdd.t28 57.8685
R62 vdd.t18 vdd.t32 57.8685
R63 vdd.t26 vdd.t30 57.8685
R64 vdd.t30 vdd.t16 57.8685
R65 vdd.t16 vdd.t22 57.8685
R66 vdd.t22 vdd.t14 57.8685
R67 vdd.t4 vdd.t43 57.8685
R68 vdd.t41 vdd.t4 57.8685
R69 vdd.t6 vdd.t41 57.8685
R70 vdd.t8 vdd.t6 57.8685
R71 vdd.t0 vdd.t2 57.8685
R72 vdd.t12 vdd.t0 57.8685
R73 vdd.t37 vdd.t12 57.8685
R74 vdd.t39 vdd.t37 57.8685
R75 vdd.n5 vdd.n3 43.602
R76 vdd.n18 vdd.n16 43.6015
R77 vdd.n23 vdd.n15 43.5947
R78 vdd.n10 vdd.n2 42.9666
R79 vdd.n18 vdd.n17 42.9638
R80 vdd.n9 vdd.n8 42.9638
R81 vdd.n20 vdd.n19 42.9611
R82 vdd.n7 vdd.n6 42.9611
R83 vdd.n22 vdd.n21 42.9584
R84 vdd.n5 vdd.n4 42.9584
R85 vdd.n14 vdd.t18 28.9345
R86 vdd.n14 vdd.t26 28.9345
R87 vdd.n11 vdd.t8 28.9345
R88 vdd.t2 vdd.n11 28.9345
R89 vdd vdd.n14 24.6672
R90 vdd.n11 vdd 24.6672
R91 vdd.n26 vdd.n25 16.0919
R92 vdd.n12 vdd.n1 16.0005
R93 vdd.n24 vdd.n23 14.8702
R94 vdd.n21 vdd.t29 5.71315
R95 vdd.n21 vdd.t33 5.71315
R96 vdd.n19 vdd.t19 5.71315
R97 vdd.n19 vdd.t27 5.71315
R98 vdd.n17 vdd.t31 5.71315
R99 vdd.n17 vdd.t17 5.71315
R100 vdd.n16 vdd.t23 5.71315
R101 vdd.n16 vdd.t15 5.71315
R102 vdd.n15 vdd.t25 5.71315
R103 vdd.n15 vdd.t21 5.71315
R104 vdd.n2 vdd.t44 5.71315
R105 vdd.n2 vdd.t5 5.71315
R106 vdd.n8 vdd.t42 5.71315
R107 vdd.n8 vdd.t7 5.71315
R108 vdd.n6 vdd.t9 5.71315
R109 vdd.n6 vdd.t3 5.71315
R110 vdd.n4 vdd.t1 5.71315
R111 vdd.n4 vdd.t13 5.71315
R112 vdd.n3 vdd.t38 5.71315
R113 vdd.n3 vdd.t40 5.71315
R114 vdd.n13 vdd 1.8768
R115 vdd.n0 vdd 1.8768
R116 vdd vdd.n26 0.731929
R117 vdd vdd.n12 0.711611
R118 vdd.n20 vdd.n18 0.64677
R119 vdd.n9 vdd.n7 0.64677
R120 vdd.n10 vdd.n9 0.625937
R121 vdd.n22 vdd 0.42212
R122 vdd vdd.n5 0.42212
R123 vdd vdd.n20 0.209999
R124 vdd.n7 vdd 0.209999
R125 vdd.n23 vdd.n22 0.00771154
R126 gnd.n21 gnd.t12 21204.1
R127 gnd.t15 gnd.n10 2972.68
R128 gnd.n19 gnd.t13 2972.68
R129 gnd.n3 gnd.t2 2340.43
R130 gnd.n18 gnd.n1 1582.12
R131 gnd.n3 gnd.t12 941.371
R132 gnd.n22 gnd.t2 748.937
R133 gnd.n9 gnd.n7 610.077
R134 gnd.n21 gnd.t6 591.941
R135 gnd.n3 gnd 585
R136 gnd gnd.n3 585
R137 gnd gnd.n22 585
R138 gnd.n21 gnd.t15 271.091
R139 gnd.n21 gnd.t13 271.091
R140 gnd.n20 gnd.n16 262.457
R141 gnd.t6 gnd.t0 261.873
R142 gnd.t0 gnd.t4 261.873
R143 gnd.t4 gnd.t8 261.873
R144 gnd.t8 gnd.t10 261.873
R145 gnd.n5 gnd.n1 237.554
R146 gnd.n2 gnd.t3 220.511
R147 gnd.t4 gnd 149.262
R148 gnd.n4 gnd 141.554
R149 gnd gnd.n20 125.919
R150 gnd.n18 gnd.n17 86.2123
R151 gnd.n9 gnd.n8 85.4593
R152 gnd.n10 gnd.n9 79.3187
R153 gnd.n5 gnd.n4 79.0593
R154 gnd.n19 gnd.n18 75.9301
R155 gnd.n20 gnd 67.9339
R156 gnd.n6 gnd.n5 61.7417
R157 gnd.n17 gnd.t14 59.2356
R158 gnd.n8 gnd.t16 59.2356
R159 gnd gnd.n1 57.7834
R160 gnd.n7 gnd.n0 57.0519
R161 gnd.n22 gnd.n21 46.809
R162 gnd.n7 gnd.n6 44.0476
R163 gnd.n6 gnd.n2 42.9181
R164 gnd.n0 gnd 33.1299
R165 gnd.n4 gnd 17.3181
R166 gnd.n15 gnd.n14 17.2621
R167 gnd.n13 gnd.n12 17.2594
R168 gnd.n16 gnd.t7 14.2966
R169 gnd.n2 gnd 9.30322
R170 gnd.n16 gnd.n15 6.98618
R171 gnd.n14 gnd.t1 3.41429
R172 gnd.n14 gnd.t5 3.41429
R173 gnd.n12 gnd.t9 3.41429
R174 gnd.n12 gnd.t11 3.41429
R175 gnd.n17 gnd 3.11409
R176 gnd.n8 gnd 3.11409
R177 gnd gnd.n0 0.731929
R178 gnd.n15 gnd.n13 0.602263
R179 gnd.n11 gnd 0.532643
R180 gnd.n10 gnd 0.420172
R181 gnd gnd.n19 0.366214
R182 gnd.n11 gnd 0.358673
R183 gnd.n13 gnd.n11 0.0774231
R184 X.n0 X.t8 1150.05
R185 X.n8 X.t3 1149.4
R186 X.n7 X.t5 1149.4
R187 X.n6 X.t9 1149.4
R188 X.n5 X.t2 1149.4
R189 X.n4 X.t7 1149.4
R190 X.n3 X.t4 1149.4
R191 X.n2 X.t10 1149.4
R192 X.n1 X.t6 1149.4
R193 X.n0 X.t11 1149.4
R194 X X.t1 117.391
R195 X.n10 X.t0 111.635
R196 X.n4 X.n3 6.02208
R197 X.n9 X 1.88686
R198 X X.n8 1.86285
R199 X.n10 X.n9 0.750006
R200 X.n1 X.n0 0.650756
R201 X.n2 X.n1 0.650756
R202 X.n3 X.n2 0.650756
R203 X.n5 X.n4 0.650756
R204 X.n7 X.n6 0.650756
R205 X.n9 X 0.637522
R206 X.n8 X.n7 0.626312
R207 X X.n5 0.340334
R208 X.n6 X 0.310922
R209 X X.n10 0.00593478
R210 vout2 vout2.t10 62.3383
R211 vout2.n1 vout2.t7 44.8719
R212 vout2.n6 vout2.t8 42.8569
R213 vout2.n1 vout2.n0 38.6225
R214 vout2.n3 vout2.n2 38.6225
R215 vout2.n8 vout2.n4 38.6225
R216 vout2.n7 vout2.n5 38.6225
R217 vout2.n0 vout2.t4 5.71315
R218 vout2.n0 vout2.t1 5.71315
R219 vout2.n2 vout2.t9 5.71315
R220 vout2.n2 vout2.t5 5.71315
R221 vout2.n4 vout2.t2 5.71315
R222 vout2.n4 vout2.t0 5.71315
R223 vout2.n5 vout2.t6 5.71315
R224 vout2.n5 vout2.t3 5.71315
R225 vout2.n7 vout2.n6 2.01553
R226 vout2.n6 vout2 1.62369
R227 vout2.n3 vout2.n1 0.537265
R228 vout2.n8 vout2.n7 0.537265
R229 vout2 vout2.n3 0.276235
R230 vout2 vout2.n8 0.261529
R231 vin1.n0 vin1.t0 358.921
R232 vin1.n0 vin1 0.0673103
R233 vin1 vin1.n0 0.00481034
R234 vin2 vin2.t0 358.925
R235 vb1 vb1.t0 599.926
R236 vb1 vb1.t1 599.926
R237 vb2.n0 vb2.t1 436.041
R238 vb2.n1 vb2.t0 436.041
R239 vb2 vb2.n0 2.91443
R240 vb2.n1 vb2 2.19389
R241 vb2 vb2.n1 0.0113696
R242 vb2.n0 vb2 0.0111383
C0 X vb1 0.09222f
C1 X vdd 2.33915f
C2 vout2 vin2 0
C3 vout1 sky130_fd_pr__nfet_01v8_DAKYLM_1.D 0.91919f
C4 vin1 Y 0.02986f
C5 vin1 vb2 0
C6 sky130_fd_pr__nfet_01v8_5Y6VJK_0.D sky130_fd_pr__nfet_01v8_DAKYLM_1.D 0.12898f
C7 vb1 vout1 0.00121f
C8 vin2 vb2 0.00198f
C9 vin2 Y 0
C10 vdd vout1 8.15727f
C11 X vin1 0
C12 vb1 sky130_fd_pr__nfet_01v8_5Y6VJK_0.D 0.06616f
C13 vb1 sky130_fd_pr__nfet_01v8_DAKYLM_1.D 0.17637f
C14 vout2 vb2 0.03453f
C15 sky130_fd_pr__nfet_01v8_5Y6VJK_0.D vdd 0.0283f
C16 vdd sky130_fd_pr__nfet_01v8_DAKYLM_1.D 0.69845f
C17 X vin2 0.03309f
C18 vb1 vdd 0.32417f
C19 vout2 X 1.41382f
C20 Y vb2 0.00118f
C21 vin1 vout1 0
C22 vin1 sky130_fd_pr__nfet_01v8_5Y6VJK_0.D 0.01494f
C23 vin1 sky130_fd_pr__nfet_01v8_DAKYLM_1.D 0
C24 X vb2 0
C25 X Y 0.01899f
C26 vin2 sky130_fd_pr__nfet_01v8_5Y6VJK_0.D 0.01498f
C27 vout2 vout1 0
C28 vb1 vin1 0.00681f
C29 vin1 vdd 0.0201f
C30 vb1 vin2 0.003f
C31 vout2 sky130_fd_pr__nfet_01v8_5Y6VJK_0.D 0.01051f
C32 vout2 sky130_fd_pr__nfet_01v8_DAKYLM_1.D 0.00303f
C33 vin2 vdd 0.02162f
C34 vout2 vb1 0.01201f
C35 Y vout1 1.4029f
C36 vb2 vout1 0.02154f
C37 vout2 vdd 8.25189f
C38 Y sky130_fd_pr__nfet_01v8_5Y6VJK_0.D 0.13942f
C39 sky130_fd_pr__nfet_01v8_5Y6VJK_0.D vb2 0.06217f
C40 vb2 sky130_fd_pr__nfet_01v8_DAKYLM_1.D 0.10553f
C41 Y sky130_fd_pr__nfet_01v8_DAKYLM_1.D 0.44045f
C42 vb1 Y 0.09067f
C43 vb1 vb2 0.07296f
C44 vin1 vin2 0.01336f
C45 X sky130_fd_pr__nfet_01v8_5Y6VJK_0.D 0.13933f
C46 X sky130_fd_pr__nfet_01v8_DAKYLM_1.D 0
C47 vb2 vdd 0.02868f
C48 Y vdd 2.64617f
C49 vout2 gnd 1.35696f
C50 vb2 gnd 0.97794f
C51 vin2 gnd 0.16094f
C52 vin1 gnd 0.16168f
C53 vb1 gnd 0.40494f
C54 vout1 gnd 2.0423f
C55 vdd gnd 18.2685f
C56 X gnd 1.51625f
C57 sky130_fd_pr__nfet_01v8_5Y6VJK_0.D gnd 0.5547f
C58 Y gnd 1.63249f
C59 sky130_fd_pr__nfet_01v8_DAKYLM_1.D gnd 7.1698f
C60 vout2.t7 gnd 0.53263f
C61 vout2.t4 gnd 0.14676f
C62 vout2.t1 gnd 0.14676f
C63 vout2.n0 gnd 0.32132f
C64 vout2.n1 gnd 1.47653f
C65 vout2.t9 gnd 0.14676f
C66 vout2.t5 gnd 0.14676f
C67 vout2.n2 gnd 0.32132f
C68 vout2.n3 gnd 0.71522f
C69 vout2.t2 gnd 0.14676f
C70 vout2.t0 gnd 0.14676f
C71 vout2.n4 gnd 0.32132f
C72 vout2.t6 gnd 0.14676f
C73 vout2.t3 gnd 0.14676f
C74 vout2.n5 gnd 0.32132f
C75 vout2.t10 gnd 0.10616f
C76 vout2.t8 gnd 0.50163f
C77 vout2.n6 gnd 0.609f
C78 vout2.n7 gnd 0.81722f
C79 vout2.n8 gnd 0.71469f
C80 X.t8 gnd 0.09579f
C81 X.t11 gnd 0.09575f
C82 X.n0 gnd 0.13685f
C83 X.t6 gnd 0.09575f
C84 X.n1 gnd 0.07243f
C85 X.t10 gnd 0.09575f
C86 X.n2 gnd 0.07243f
C87 X.t4 gnd 0.09575f
C88 X.n3 gnd 0.16138f
C89 X.t7 gnd 0.09575f
C90 X.n4 gnd 0.16114f
C91 X.t2 gnd 0.09575f
C92 X.n5 gnd 0.06716f
C93 X.t9 gnd 0.09575f
C94 X.n6 gnd 0.06666f
C95 X.t5 gnd 0.09575f
C96 X.n7 gnd 0.0726f
C97 X.t3 gnd 0.09575f
C98 X.n8 gnd 0.09532f
C99 X.t1 gnd 0.03121f
C100 X.n9 gnd 0.0576f
C101 X.t0 gnd 0.08502f
C102 X.n10 gnd 0.10035f
C103 vdd.t11 gnd 0.07038f
C104 vdd.n0 gnd 0.04484f
C105 vdd.n1 gnd 0.06585f
C106 vdd.t43 gnd 1.21171f
C107 vdd.t4 gnd 0.4423f
C108 vdd.t41 gnd 0.4423f
C109 vdd.t6 gnd 0.4423f
C110 vdd.t8 gnd 0.33172f
C111 vdd.t44 gnd 0.05489f
C112 vdd.t5 gnd 0.05489f
C113 vdd.n2 gnd 0.14193f
C114 vdd.t38 gnd 0.05489f
C115 vdd.t40 gnd 0.05489f
C116 vdd.n3 gnd 0.14502f
C117 vdd.t1 gnd 0.05489f
C118 vdd.t13 gnd 0.05489f
C119 vdd.n4 gnd 0.14181f
C120 vdd.n5 gnd 0.43865f
C121 vdd.t9 gnd 0.05489f
C122 vdd.t3 gnd 0.05489f
C123 vdd.n6 gnd 0.14185f
C124 vdd.n7 gnd 0.21989f
C125 vdd.t42 gnd 0.05489f
C126 vdd.t7 gnd 0.05489f
C127 vdd.n8 gnd 0.14189f
C128 vdd.n9 gnd 0.22606f
C129 vdd.n10 gnd 0.29684f
C130 vdd.n11 gnd 0.48534f
C131 vdd.t2 gnd 0.33172f
C132 vdd.t0 gnd 0.4423f
C133 vdd.t12 gnd 0.4423f
C134 vdd.t37 gnd 0.4423f
C135 vdd.t39 gnd 1.1106f
C136 vdd.t10 gnd 0.92571f
C137 vdd.n12 gnd 0.39709f
C138 vdd.t35 gnd 0.07038f
C139 vdd.n13 gnd 0.04488f
C140 vdd.t36 gnd 0.1013f
C141 vdd.t24 gnd 1.21171f
C142 vdd.t20 gnd 0.4423f
C143 vdd.t28 gnd 0.4423f
C144 vdd.t32 gnd 0.4423f
C145 vdd.t18 gnd 0.33172f
C146 vdd.t14 gnd 1.21171f
C147 vdd.t22 gnd 0.4423f
C148 vdd.t16 gnd 0.4423f
C149 vdd.t30 gnd 0.4423f
C150 vdd.t26 gnd 0.33172f
C151 vdd.n14 gnd 0.48534f
C152 vdd.t25 gnd 0.05489f
C153 vdd.t21 gnd 0.05489f
C154 vdd.n15 gnd 0.14498f
C155 vdd.t23 gnd 0.05489f
C156 vdd.t15 gnd 0.05489f
C157 vdd.n16 gnd 0.14514f
C158 vdd.t31 gnd 0.05489f
C159 vdd.t17 gnd 0.05489f
C160 vdd.n17 gnd 0.14189f
C161 vdd.n18 gnd 0.4429f
C162 vdd.t19 gnd 0.05489f
C163 vdd.t27 gnd 0.05489f
C164 vdd.n19 gnd 0.14185f
C165 vdd.n20 gnd 0.21989f
C166 vdd.t29 gnd 0.05489f
C167 vdd.t33 gnd 0.05489f
C168 vdd.n21 gnd 0.14181f
C169 vdd.n22 gnd 0.21173f
C170 vdd.n23 gnd 0.26543f
C171 vdd.n24 gnd 0.09101f
C172 vdd.n25 gnd 0.09499f
C173 vdd.t34 gnd 0.8246f
C174 vdd.n26 gnd 0.39698f
C175 vout1.t3 gnd 0.13772f
C176 vout1.t8 gnd 0.13772f
C177 vout1.n0 gnd 0.30155f
C178 vout1.t2 gnd 0.13772f
C179 vout1.t5 gnd 0.13772f
C180 vout1.n1 gnd 0.30155f
C181 vout1.t10 gnd 0.09963f
C182 vout1.t9 gnd 0.47076f
C183 vout1.n2 gnd 0.60805f
C184 vout1.n3 gnd 0.76692f
C185 vout1.n4 gnd 0.67071f
C186 vout1.t6 gnd 0.49985f
C187 vout1.t4 gnd 0.13772f
C188 vout1.t7 gnd 0.13772f
C189 vout1.n5 gnd 0.30155f
C190 vout1.n6 gnd 1.38566f
C191 vout1.t1 gnd 0.13772f
C192 vout1.t0 gnd 0.13772f
C193 vout1.n7 gnd 0.30155f
C194 vout1.n8 gnd 0.6712f
C195 Y.t6 gnd 0.10284f
C196 Y.t8 gnd 0.10288f
C197 Y.t2 gnd 0.10284f
C198 Y.n0 gnd 0.14698f
C199 Y.t5 gnd 0.10284f
C200 Y.n1 gnd 0.07778f
C201 Y.t10 gnd 0.10284f
C202 Y.n2 gnd 0.07778f
C203 Y.t11 gnd 0.10284f
C204 Y.n3 gnd 0.17332f
C205 Y.t7 gnd 0.10284f
C206 Y.n4 gnd 0.17307f
C207 Y.t3 gnd 0.10284f
C208 Y.n5 gnd 0.07213f
C209 Y.t9 gnd 0.10284f
C210 Y.n6 gnd 0.0716f
C211 Y.t4 gnd 0.10284f
C212 Y.n7 gnd 0.07762f
C213 Y.n8 gnd 0.1664f
C214 Y.t1 gnd 0.03352f
C215 Y.n9 gnd 0.07274f
C216 Y.t0 gnd 0.09131f
C217 Y.n10 gnd 0.09894f
.ends

