magic
tech sky130A
magscale 1 2
timestamp 1719358519
<< nwell >>
rect -647 -788 647 788
<< pmos >>
rect -447 -569 -417 569
rect -351 -569 -321 569
rect -255 -569 -225 569
rect -159 -569 -129 569
rect -63 -569 -33 569
rect 33 -569 63 569
rect 129 -569 159 569
rect 225 -569 255 569
rect 321 -569 351 569
rect 417 -569 447 569
<< pdiff >>
rect -509 557 -447 569
rect -509 -557 -497 557
rect -463 -557 -447 557
rect -509 -569 -447 -557
rect -417 557 -351 569
rect -417 -557 -401 557
rect -367 -557 -351 557
rect -417 -569 -351 -557
rect -321 557 -255 569
rect -321 -557 -305 557
rect -271 -557 -255 557
rect -321 -569 -255 -557
rect -225 557 -159 569
rect -225 -557 -209 557
rect -175 -557 -159 557
rect -225 -569 -159 -557
rect -129 557 -63 569
rect -129 -557 -113 557
rect -79 -557 -63 557
rect -129 -569 -63 -557
rect -33 557 33 569
rect -33 -557 -17 557
rect 17 -557 33 557
rect -33 -569 33 -557
rect 63 557 129 569
rect 63 -557 79 557
rect 113 -557 129 557
rect 63 -569 129 -557
rect 159 557 225 569
rect 159 -557 175 557
rect 209 -557 225 557
rect 159 -569 225 -557
rect 255 557 321 569
rect 255 -557 271 557
rect 305 -557 321 557
rect 255 -569 321 -557
rect 351 557 417 569
rect 351 -557 367 557
rect 401 -557 417 557
rect 351 -569 417 -557
rect 447 557 509 569
rect 447 -557 463 557
rect 497 -557 509 557
rect 447 -569 509 -557
<< pdiffc >>
rect -497 -557 -463 557
rect -401 -557 -367 557
rect -305 -557 -271 557
rect -209 -557 -175 557
rect -113 -557 -79 557
rect -17 -557 17 557
rect 79 -557 113 557
rect 175 -557 209 557
rect 271 -557 305 557
rect 367 -557 401 557
rect 463 -557 497 557
<< nsubdiff >>
rect -611 718 -515 752
rect 515 718 611 752
rect -611 -718 -577 718
rect 577 -718 611 718
rect -611 -752 611 -718
<< nsubdiffcont >>
rect -515 718 515 752
<< poly >>
rect -369 650 -303 666
rect -369 616 -353 650
rect -319 616 -303 650
rect -369 600 -303 616
rect -177 650 -111 666
rect -177 616 -161 650
rect -127 616 -111 650
rect -177 600 -111 616
rect 15 650 81 666
rect 15 616 31 650
rect 65 616 81 650
rect 15 600 81 616
rect 207 650 273 666
rect 207 616 223 650
rect 257 616 273 650
rect 207 600 273 616
rect 399 650 465 666
rect 399 616 415 650
rect 449 616 465 650
rect 399 600 465 616
rect -447 569 -417 595
rect -351 569 -321 600
rect -255 569 -225 595
rect -159 569 -129 600
rect -63 569 -33 595
rect 33 569 63 600
rect 129 569 159 595
rect 225 569 255 600
rect 321 569 351 595
rect 417 569 447 600
rect -447 -600 -417 -569
rect -351 -595 -321 -569
rect -255 -600 -225 -569
rect -159 -595 -129 -569
rect -63 -600 -33 -569
rect 33 -595 63 -569
rect 129 -600 159 -569
rect 225 -595 255 -569
rect 321 -600 351 -569
rect 417 -595 447 -569
rect -465 -616 -399 -600
rect -465 -650 -449 -616
rect -415 -650 -399 -616
rect -465 -666 -399 -650
rect -273 -616 -207 -600
rect -273 -650 -257 -616
rect -223 -650 -207 -616
rect -273 -666 -207 -650
rect -81 -616 -15 -600
rect -81 -650 -65 -616
rect -31 -650 -15 -616
rect -81 -666 -15 -650
rect 111 -616 177 -600
rect 111 -650 127 -616
rect 161 -650 177 -616
rect 111 -666 177 -650
rect 303 -616 369 -600
rect 303 -650 319 -616
rect 353 -650 369 -616
rect 303 -666 369 -650
<< polycont >>
rect -353 616 -319 650
rect -161 616 -127 650
rect 31 616 65 650
rect 223 616 257 650
rect 415 616 449 650
rect -449 -650 -415 -616
rect -257 -650 -223 -616
rect -65 -650 -31 -616
rect 127 -650 161 -616
rect 319 -650 353 -616
<< locali >>
rect -531 718 -515 752
rect 515 718 531 752
rect -369 616 -353 650
rect -319 616 -303 650
rect -177 616 -161 650
rect -127 616 -111 650
rect 15 616 31 650
rect 65 616 81 650
rect 207 616 223 650
rect 257 616 273 650
rect 399 616 415 650
rect 449 616 465 650
rect -497 557 -463 573
rect -497 -573 -463 -557
rect -401 557 -367 573
rect -401 -573 -367 -557
rect -305 557 -271 573
rect -305 -573 -271 -557
rect -209 557 -175 573
rect -209 -573 -175 -557
rect -113 557 -79 573
rect -113 -573 -79 -557
rect -17 557 17 573
rect -17 -573 17 -557
rect 79 557 113 573
rect 79 -573 113 -557
rect 175 557 209 573
rect 175 -573 209 -557
rect 271 557 305 573
rect 271 -573 305 -557
rect 367 557 401 573
rect 367 -573 401 -557
rect 463 557 497 573
rect 463 -573 497 -557
rect -465 -650 -449 -616
rect -415 -650 -399 -616
rect -273 -650 -257 -616
rect -223 -650 -207 -616
rect -81 -650 -65 -616
rect -31 -650 -15 -616
rect 111 -650 127 -616
rect 161 -650 177 -616
rect 303 -650 319 -616
rect 353 -650 369 -616
<< viali >>
rect -353 616 -319 650
rect -161 616 -127 650
rect 31 616 65 650
rect 223 616 257 650
rect 415 616 449 650
rect -497 -557 -463 557
rect -401 -446 -367 446
rect -305 -557 -271 557
rect -209 -446 -175 446
rect -113 -557 -79 557
rect -17 -446 17 446
rect 79 -557 113 557
rect 175 -446 209 446
rect 271 -557 305 557
rect 367 -446 401 446
rect 463 -557 497 557
rect -449 -650 -415 -616
rect -257 -650 -223 -616
rect -65 -650 -31 -616
rect 127 -650 161 -616
rect 319 -650 353 -616
<< metal1 >>
rect -365 653 -307 656
rect -173 653 -115 656
rect 19 653 77 656
rect 211 653 269 656
rect 403 653 461 656
rect -610 650 461 653
rect -610 619 -353 650
rect -610 -616 -576 619
rect -365 616 -353 619
rect -319 619 -161 650
rect -319 616 -307 619
rect -365 610 -307 616
rect -173 616 -161 619
rect -127 619 31 650
rect -127 616 -115 619
rect -173 610 -115 616
rect 19 616 31 619
rect 65 619 223 650
rect 65 616 77 619
rect 19 610 77 616
rect 211 616 223 619
rect 257 619 415 650
rect 257 616 269 619
rect 211 610 269 616
rect 403 616 415 619
rect 449 616 461 650
rect 403 610 461 616
rect -503 561 -457 569
rect -311 561 -265 569
rect -119 561 -73 569
rect 73 561 119 569
rect 265 561 311 569
rect 457 561 503 569
rect -503 557 503 561
rect -503 -557 -497 557
rect -463 527 -305 557
rect -463 -557 -457 527
rect -407 451 -361 458
rect -410 446 -358 451
rect -410 445 -401 446
rect -367 445 -358 446
rect -410 387 -401 393
rect -407 -446 -401 387
rect -367 387 -358 393
rect -367 -446 -361 387
rect -407 -458 -361 -446
rect -503 -569 -457 -557
rect -311 -557 -305 527
rect -271 527 -113 557
rect -271 -557 -265 527
rect -215 450 -169 458
rect -219 446 -167 450
rect -219 444 -209 446
rect -175 444 -167 446
rect -219 386 -209 392
rect -215 -446 -209 386
rect -175 386 -167 392
rect -175 -446 -169 386
rect -215 -458 -169 -446
rect -311 -569 -265 -557
rect -119 -557 -113 527
rect -79 527 79 557
rect -79 -557 -73 527
rect -23 449 23 458
rect -25 446 27 449
rect -25 443 -17 446
rect 17 443 27 446
rect -25 385 -17 391
rect -23 -446 -17 385
rect 17 385 27 391
rect 17 -446 23 385
rect -23 -458 23 -446
rect -119 -569 -73 -557
rect 73 -557 79 527
rect 113 527 271 557
rect 113 -557 119 527
rect 169 448 215 458
rect 165 446 217 448
rect 165 442 175 446
rect 209 442 217 446
rect 165 384 175 390
rect 169 -446 175 384
rect 209 384 217 390
rect 209 -446 215 384
rect 169 -458 215 -446
rect 73 -569 119 -557
rect 265 -557 271 527
rect 305 527 463 557
rect 305 -557 311 527
rect 361 447 407 458
rect 359 446 411 447
rect 359 441 367 446
rect 401 441 411 446
rect 359 383 367 389
rect 361 -446 367 383
rect 401 383 411 389
rect 401 -446 407 383
rect 361 -458 407 -446
rect 265 -569 311 -557
rect 457 -557 463 527
rect 497 -557 503 557
rect 457 -569 503 -557
rect -461 -616 -403 -610
rect -269 -616 -211 -610
rect -77 -616 -19 -610
rect 115 -616 173 -610
rect 307 -616 365 -610
rect -610 -650 -449 -616
rect -415 -650 -257 -616
rect -223 -650 -65 -616
rect -31 -650 127 -616
rect 161 -650 319 -616
rect 353 -650 365 -616
rect -461 -656 -403 -650
rect -269 -656 -211 -650
rect -77 -656 -19 -650
rect 115 -656 173 -650
rect 307 -656 365 -650
<< via1 >>
rect -410 393 -401 445
rect -401 393 -367 445
rect -367 393 -358 445
rect -219 392 -209 444
rect -209 392 -175 444
rect -175 392 -167 444
rect -25 391 -17 443
rect -17 391 17 443
rect 17 391 27 443
rect 165 390 175 442
rect 175 390 209 442
rect 209 390 217 442
rect 359 389 367 441
rect 367 389 401 441
rect 401 389 411 441
<< metal2 >>
rect -416 393 -410 445
rect -358 435 -352 445
rect -225 435 -219 444
rect -358 402 -219 435
rect -358 393 -352 402
rect -225 392 -219 402
rect -167 434 -161 444
rect -31 434 -25 443
rect -167 401 -25 434
rect -167 392 -161 401
rect -31 391 -25 401
rect 27 433 33 443
rect 159 433 165 442
rect 27 400 165 433
rect 27 391 33 400
rect 159 390 165 400
rect 217 432 223 442
rect 353 432 359 441
rect 217 399 359 432
rect 217 390 223 399
rect 353 389 359 399
rect 411 389 417 441
<< labels >>
flabel metal1 s 2 549 2 549 0 FreeSans 480 0 0 0 D
port 0 nsew
flabel metal2 s 68 416 68 416 0 FreeSans 480 0 0 0 S
port 1 nsew
flabel metal1 s -44 632 -44 632 0 FreeSans 480 0 0 0 G
port 2 nsew
flabel locali s 0 736 0 736 0 FreeSans 480 0 0 0 B
port 3 nsew
<< properties >>
string FIXED_BBOX -594 -735 594 735
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 5.69 l 0.15 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 1 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 80 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
