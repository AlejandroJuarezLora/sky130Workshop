* NGSPICE file created from opamp.ext - technology: sky130B

.subckt opamp_pex vdd gnd vout2 vout1 vb2 vb1 vin1 vin2
X0 vdd.t21 Y.t2 vout1.t0 vdd.t20 sky130_fd_pr__pfet_01v8 ad=0.93885 pd=6.02 as=0.93885 ps=6.02 w=5.69 l=0.15
X1 gnd.t11 sky130_fd_pr__nfet_01v8_DAKYLM_1.D sky130_fd_pr__nfet_01v8_DAKYLM_1.D gnd.t10 sky130_fd_pr__nfet_01v8 ad=0.957 pd=6.13 as=1.798 ps=12.22 w=5.8 l=0.15
X2 gnd.t9 sky130_fd_pr__nfet_01v8_DAKYLM_1.D sky130_fd_pr__nfet_01v8_5Y6VJK_0.D gnd.t8 sky130_fd_pr__nfet_01v8 ad=0.1421 pd=1.56 as=0.1421 ps=1.56 w=0.49 l=0.15
X3 vout1.t1 Y.t3 vdd.t19 vdd.t18 sky130_fd_pr__pfet_01v8 ad=0.93885 pd=6.02 as=0.93885 ps=6.02 w=5.69 l=0.15
X4 vdd.t43 X.t2 vout2.t10 vdd.t42 sky130_fd_pr__pfet_01v8 ad=0.93885 pd=6.02 as=0.93885 ps=6.02 w=5.69 l=0.15
X5 vdd.t41 X.t3 vout2.t9 vdd.t40 sky130_fd_pr__pfet_01v8 ad=0.93885 pd=6.02 as=1.7639 ps=12 w=5.69 l=0.15
X6 vout1.t4 Y.t4 vdd.t17 vdd.t16 sky130_fd_pr__pfet_01v8 ad=0.93885 pd=6.02 as=0.93885 ps=6.02 w=5.69 l=0.15
X7 sky130_fd_pr__nfet_01v8_DAKYLM_1.D sky130_fd_pr__nfet_01v8_DAKYLM_1.D gnd.t7 gnd.t6 sky130_fd_pr__nfet_01v8 ad=0.957 pd=6.13 as=0.957 ps=6.13 w=5.8 l=0.15
X8 sky130_fd_pr__nfet_01v8_5Y6VJK_0.D vin1.t0 Y.t0 gnd.t12 sky130_fd_pr__nfet_01v8 ad=0.2494 pd=2.3 as=0.2494 ps=2.3 w=0.86 l=0.15
X9 X.t1 vin2.t0 sky130_fd_pr__nfet_01v8_5Y6VJK_0.D gnd.t12 sky130_fd_pr__nfet_01v8 ad=0.2494 pd=2.3 as=0.2494 ps=2.3 w=0.86 l=0.15
X10 vdd.t15 Y.t5 vout1.t8 vdd.t14 sky130_fd_pr__pfet_01v8 ad=0.93885 pd=6.02 as=0.93885 ps=6.02 w=5.69 l=0.15
X11 vout1.t2 Y.t6 vdd.t13 vdd.t12 sky130_fd_pr__pfet_01v8 ad=1.7639 pd=12 as=0.93885 ps=6.02 w=5.69 l=0.15
X12 Y.t1 vb1.t0 vdd.t23 vdd.t22 sky130_fd_pr__pfet_01v8 ad=0.6583 pd=5.12 as=0.6583 ps=5.12 w=2.27 l=0.15
X13 vout1.t7 Y.t7 vdd.t11 vdd.t10 sky130_fd_pr__pfet_01v8 ad=0.93885 pd=6.02 as=0.93885 ps=6.02 w=5.69 l=0.15
X14 gnd.t5 sky130_fd_pr__nfet_01v8_DAKYLM_1.D sky130_fd_pr__nfet_01v8_DAKYLM_1.D gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.798 pd=12.22 as=0.957 ps=6.13 w=5.8 l=0.15
X15 vout2.t8 X.t4 vdd.t39 vdd.t38 sky130_fd_pr__pfet_01v8 ad=1.7639 pd=12 as=0.93885 ps=6.02 w=5.69 l=0.15
R0 vdd sky130_fd_pr__nfet_01v8_DAKYLM_1.D sky130_fd_pr__res_generic_po w=0.33 l=1.65
X16 vdd.t9 Y.t8 vout1.t6 vdd.t8 sky130_fd_pr__pfet_01v8 ad=0.93885 pd=6.02 as=0.93885 ps=6.02 w=5.69 l=0.15
X17 vdd.t37 X.t5 vout2.t7 vdd.t36 sky130_fd_pr__pfet_01v8 ad=0.93885 pd=6.02 as=0.93885 ps=6.02 w=5.69 l=0.15
X18 vout1.t9 Y.t9 vdd.t7 vdd.t6 sky130_fd_pr__pfet_01v8 ad=0.93885 pd=6.02 as=0.93885 ps=6.02 w=5.69 l=0.15
X19 vout2.t6 X.t6 vdd.t35 vdd.t34 sky130_fd_pr__pfet_01v8 ad=0.93885 pd=6.02 as=0.93885 ps=6.02 w=5.69 l=0.15
X20 vdd.t5 Y.t10 vout1.t3 vdd.t4 sky130_fd_pr__pfet_01v8 ad=0.93885 pd=6.02 as=0.93885 ps=6.02 w=5.69 l=0.15
X21 vdd.t1 vb1.t1 X.t0 vdd.t0 sky130_fd_pr__pfet_01v8 ad=0.6583 pd=5.12 as=0.6583 ps=5.12 w=2.27 l=0.15
X22 vdd.t33 X.t7 vout2.t5 vdd.t32 sky130_fd_pr__pfet_01v8 ad=0.93885 pd=6.02 as=0.93885 ps=6.02 w=5.69 l=0.15
X23 vout2.t4 X.t8 vdd.t31 vdd.t30 sky130_fd_pr__pfet_01v8 ad=0.93885 pd=6.02 as=0.93885 ps=6.02 w=5.69 l=0.15
X24 gnd.t3 sky130_fd_pr__nfet_01v8_DAKYLM_1.D sky130_fd_pr__nfet_01v8_DAKYLM_1.D gnd.t2 sky130_fd_pr__nfet_01v8 ad=0.957 pd=6.13 as=0.957 ps=6.13 w=5.8 l=0.15
X25 gnd.t16 vb2.t0 vout1.t10 gnd.t15 sky130_fd_pr__nfet_01v8 ad=0.3886 pd=3.26 as=0.3886 ps=3.26 w=1.34 l=0.15
X26 vdd.t29 X.t9 vout2.t3 vdd.t28 sky130_fd_pr__pfet_01v8 ad=0.93885 pd=6.02 as=0.93885 ps=6.02 w=5.69 l=0.15
X27 vout2.t0 vb2.t1 gnd.t14 gnd.t13 sky130_fd_pr__nfet_01v8 ad=0.3886 pd=3.26 as=0.3886 ps=3.26 w=1.34 l=0.15
X28 vout2.t2 X.t10 vdd.t27 vdd.t26 sky130_fd_pr__pfet_01v8 ad=0.93885 pd=6.02 as=0.93885 ps=6.02 w=5.69 l=0.15
X29 vdd.t3 Y.t11 vout1.t5 vdd.t2 sky130_fd_pr__pfet_01v8 ad=0.93885 pd=6.02 as=1.7639 ps=12 w=5.69 l=0.15
X30 sky130_fd_pr__nfet_01v8_DAKYLM_1.D sky130_fd_pr__nfet_01v8_DAKYLM_1.D gnd.t1 gnd.t0 sky130_fd_pr__nfet_01v8 ad=0.957 pd=6.13 as=0.957 ps=6.13 w=5.8 l=0.15
X31 vout2.t1 X.t11 vdd.t25 vdd.t24 sky130_fd_pr__pfet_01v8 ad=0.93885 pd=6.02 as=0.93885 ps=6.02 w=5.69 l=0.15
R1 Y.n0 Y.t8 1150.05
R2 Y.n4 Y.t6 1149.41
R3 Y.n4 Y.t4 1149.4
R4 Y.n3 Y.t9 1149.4
R5 Y.n2 Y.t3 1149.4
R6 Y.n2 Y.t7 1149.4
R7 Y.n1 Y.t11 1149.4
R8 Y.n1 Y.t10 1149.4
R9 Y.n0 Y.t5 1149.4
R10 Y.n0 Y.t2 1149.4
R11 Y Y.t0 117.392
R12 Y Y.t1 111.635
R13 Y.n2 Y.n1 6.02208
R14 Y Y.n4 4.35576
R15 Y.n1 Y.n0 1.95127
R16 Y.n3 Y.n2 1.30101
R17 Y.n4 Y.n3 1.29286
R18 vout1 vout1.t10 62.3383
R19 vout1.n6 vout1.t5 44.8719
R20 vout1.n2 vout1.t2 42.8569
R21 vout1.n6 vout1.n5 38.6225
R22 vout1.n8 vout1.n7 38.6225
R23 vout1.n4 vout1.n0 38.6225
R24 vout1.n3 vout1.n1 38.6225
R25 vout1.n5 vout1.t3 5.71315
R26 vout1.n5 vout1.t7 5.71315
R27 vout1.n7 vout1.t8 5.71315
R28 vout1.n7 vout1.t1 5.71315
R29 vout1.n0 vout1.t0 5.71315
R30 vout1.n0 vout1.t9 5.71315
R31 vout1.n1 vout1.t6 5.71315
R32 vout1.n1 vout1.t4 5.71315
R33 vout1.n2 vout1 2.42124
R34 vout1.n3 vout1.n2 2.01553
R35 vout1.n8 vout1.n6 0.537265
R36 vout1.n4 vout1.n3 0.537265
R37 vout1 vout1.n8 0.276235
R38 vout1 vout1.n4 0.261529
R39 vdd.n26 vdd.t22 909.881
R40 vdd.n12 vdd.t0 909.881
R41 vdd.n25 vdd.n24 525.279
R42 vdd vdd.n1 324.118
R43 vdd.t0 vdd.t40 210.643
R44 vdd vdd.n10 162.881
R45 vdd.n25 vdd.n13 113.942
R46 vdd.n1 vdd.n0 112.733
R47 vdd.n13 vdd.t23 110.085
R48 vdd.n0 vdd.t1 110.085
R49 vdd.n24 vdd 74.1861
R50 vdd.t8 vdd.t12 57.8685
R51 vdd.t16 vdd.t8 57.8685
R52 vdd.t20 vdd.t16 57.8685
R53 vdd.t6 vdd.t20 57.8685
R54 vdd.t14 vdd.t18 57.8685
R55 vdd.t18 vdd.t4 57.8685
R56 vdd.t4 vdd.t10 57.8685
R57 vdd.t10 vdd.t2 57.8685
R58 vdd.t32 vdd.t38 57.8685
R59 vdd.t26 vdd.t32 57.8685
R60 vdd.t42 vdd.t26 57.8685
R61 vdd.t34 vdd.t42 57.8685
R62 vdd.t24 vdd.t28 57.8685
R63 vdd.t36 vdd.t24 57.8685
R64 vdd.t30 vdd.t36 57.8685
R65 vdd.t40 vdd.t30 57.8685
R66 vdd.n5 vdd.n3 48.102
R67 vdd.n18 vdd.n16 48.1015
R68 vdd.n23 vdd.n15 48.0947
R69 vdd.n10 vdd.n2 47.4666
R70 vdd.n18 vdd.n17 47.4638
R71 vdd.n9 vdd.n8 47.4638
R72 vdd.n20 vdd.n19 47.4611
R73 vdd.n7 vdd.n6 47.4611
R74 vdd.n22 vdd.n21 47.4584
R75 vdd.n5 vdd.n4 47.4584
R76 vdd.n14 vdd.t6 28.9345
R77 vdd.n14 vdd.t14 28.9345
R78 vdd.n11 vdd.t34 28.9345
R79 vdd.t28 vdd.n11 28.9345
R80 vdd vdd.n14 24.6672
R81 vdd.n11 vdd 24.6672
R82 vdd.n24 vdd.n23 19.3702
R83 vdd.n26 vdd.n25 16.0919
R84 vdd.n12 vdd.n1 16.0005
R85 vdd.n21 vdd.t17 5.71315
R86 vdd.n21 vdd.t21 5.71315
R87 vdd.n19 vdd.t7 5.71315
R88 vdd.n19 vdd.t15 5.71315
R89 vdd.n17 vdd.t19 5.71315
R90 vdd.n17 vdd.t5 5.71315
R91 vdd.n16 vdd.t11 5.71315
R92 vdd.n16 vdd.t3 5.71315
R93 vdd.n15 vdd.t13 5.71315
R94 vdd.n15 vdd.t9 5.71315
R95 vdd.n2 vdd.t39 5.71315
R96 vdd.n2 vdd.t33 5.71315
R97 vdd.n8 vdd.t27 5.71315
R98 vdd.n8 vdd.t43 5.71315
R99 vdd.n6 vdd.t35 5.71315
R100 vdd.n6 vdd.t29 5.71315
R101 vdd.n4 vdd.t25 5.71315
R102 vdd.n4 vdd.t37 5.71315
R103 vdd.n3 vdd.t31 5.71315
R104 vdd.n3 vdd.t41 5.71315
R105 vdd.n13 vdd 1.8768
R106 vdd.n0 vdd 1.8768
R107 vdd vdd.n26 0.731929
R108 vdd vdd.n12 0.711611
R109 vdd.n20 vdd.n18 0.64677
R110 vdd.n9 vdd.n7 0.64677
R111 vdd.n10 vdd.n9 0.625937
R112 vdd.n22 vdd 0.42212
R113 vdd vdd.n5 0.42212
R114 vdd vdd.n20 0.209999
R115 vdd.n7 vdd 0.209999
R116 vdd.n23 vdd.n22 0.00771154
R117 gnd.n21 gnd.t12 21204.1
R118 gnd.t13 gnd.n10 2972.68
R119 gnd.n19 gnd.t15 2972.68
R120 gnd.n3 gnd.t8 2340.43
R121 gnd.n18 gnd.n1 1582.12
R122 gnd.n3 gnd.t12 941.371
R123 gnd.n22 gnd.t8 748.937
R124 gnd.n9 gnd.n7 610.077
R125 gnd.n21 gnd.t4 591.941
R126 gnd.n3 gnd 585
R127 gnd gnd.n3 585
R128 gnd gnd.n22 585
R129 gnd.n21 gnd.t13 271.091
R130 gnd.n21 gnd.t15 271.091
R131 gnd.n20 gnd.n16 262.457
R132 gnd.t4 gnd.t0 261.873
R133 gnd.t0 gnd.t2 261.873
R134 gnd.t2 gnd.t6 261.873
R135 gnd.t6 gnd.t10 261.873
R136 gnd.n5 gnd.n1 237.554
R137 gnd.n2 gnd.t9 220.511
R138 gnd.t2 gnd 149.262
R139 gnd.n4 gnd 141.554
R140 gnd gnd.n20 125.919
R141 gnd.n18 gnd.n17 86.2123
R142 gnd.n9 gnd.n8 85.4593
R143 gnd.n10 gnd.n9 79.3187
R144 gnd.n5 gnd.n4 79.0593
R145 gnd.n19 gnd.n18 75.9301
R146 gnd.n20 gnd 67.9339
R147 gnd.n6 gnd.n5 61.7417
R148 gnd.n17 gnd.t16 59.2356
R149 gnd.n8 gnd.t14 59.2356
R150 gnd gnd.n1 57.7834
R151 gnd.n7 gnd.n0 57.0519
R152 gnd.n22 gnd.n21 46.809
R153 gnd.n7 gnd.n6 44.0476
R154 gnd.n6 gnd.n2 42.9181
R155 gnd.n0 gnd 33.1299
R156 gnd.n15 gnd.n14 21.7621
R157 gnd.n13 gnd.n12 21.7594
R158 gnd.n4 gnd 17.3181
R159 gnd.n16 gnd.t5 14.2966
R160 gnd.n16 gnd.n15 11.4862
R161 gnd.n2 gnd 9.30322
R162 gnd.n14 gnd.t1 3.41429
R163 gnd.n14 gnd.t3 3.41429
R164 gnd.n12 gnd.t7 3.41429
R165 gnd.n12 gnd.t11 3.41429
R166 gnd.n17 gnd 3.11409
R167 gnd.n8 gnd 3.11409
R168 gnd gnd.n0 0.731929
R169 gnd.n15 gnd.n13 0.602263
R170 gnd.n11 gnd 0.532643
R171 gnd.n10 gnd 0.420172
R172 gnd gnd.n19 0.366214
R173 gnd.n11 gnd 0.358673
R174 gnd.n13 gnd.n11 0.0774231
R175 X.n0 X.t8 1150.05
R176 X.n4 X.t3 1149.4
R177 X.n4 X.t5 1149.4
R178 X.n3 X.t9 1149.4
R179 X.n2 X.t2 1149.4
R180 X.n2 X.t7 1149.4
R181 X.n1 X.t4 1149.4
R182 X.n1 X.t10 1149.4
R183 X.n0 X.t6 1149.4
R184 X.n0 X.t11 1149.4
R185 X X.t1 117.391
R186 X X.t0 111.635
R187 X.n2 X.n1 6.02208
R188 X.n1 X.n0 1.95127
R189 X X.n4 1.86285
R190 X.n3 X.n2 1.30101
R191 X.n4 X.n3 1.27657
R192 vout2 vout2.t0 62.3383
R193 vout2.n1 vout2.t8 44.8719
R194 vout2.n6 vout2.t9 42.8569
R195 vout2.n1 vout2.n0 38.6225
R196 vout2.n3 vout2.n2 38.6225
R197 vout2.n8 vout2.n4 38.6225
R198 vout2.n7 vout2.n5 38.6225
R199 vout2.n0 vout2.t5 5.71315
R200 vout2.n0 vout2.t2 5.71315
R201 vout2.n2 vout2.t10 5.71315
R202 vout2.n2 vout2.t6 5.71315
R203 vout2.n4 vout2.t3 5.71315
R204 vout2.n4 vout2.t1 5.71315
R205 vout2.n5 vout2.t7 5.71315
R206 vout2.n5 vout2.t4 5.71315
R207 vout2.n7 vout2.n6 2.01553
R208 vout2.n6 vout2 1.62369
R209 vout2.n3 vout2.n1 0.537265
R210 vout2.n8 vout2.n7 0.537265
R211 vout2 vout2.n3 0.276235
R212 vout2 vout2.n8 0.261529
R213 vin1.n0 vin1.t0 358.921
R214 vin1.n0 vin1 0.0673103
R215 vin1 vin1.n0 0.00481034
R216 vin2 vin2.t0 358.925
R217 vb1 vb1.t0 599.926
R218 vb1 vb1.t1 599.926
R219 vb2.n0 vb2.t1 436.041
R220 vb2.n1 vb2.t0 436.041
R221 vb2 vb2.n0 2.91443
R222 vb2.n1 vb2 2.19389
R223 vb2 vb2.n1 0.0113696
R224 vb2.n0 vb2 0.0111383
C0 vout2 vin2 2.13e-19
C1 X vin1 2.23e-19
C2 sky130_fd_pr__nfet_01v8_5Y6VJK_0.D sky130_fd_pr__nfet_01v8_DAKYLM_1.D 0.093021f
C3 vb1 X 0.092133f
C4 vb2 sky130_fd_pr__nfet_01v8_DAKYLM_1.D 0.104891f
C5 sky130_fd_pr__nfet_01v8_5Y6VJK_0.D vin1 0.014938f
C6 sky130_fd_pr__nfet_01v8_5Y6VJK_0.D vb1 0.042727f
C7 vb2 vin1 5.22e-21
C8 vout2 sky130_fd_pr__nfet_01v8_DAKYLM_1.D 0.003021f
C9 Y vdd 2.60583f
C10 vb2 vout1 0.021544f
C11 vb2 vb1 0.072899f
C12 vout2 vout1 7.95e-19
C13 vout2 vb1 0.011987f
C14 X Y 0.018987f
C15 X vdd 2.29926f
C16 sky130_fd_pr__nfet_01v8_5Y6VJK_0.D Y 0.139423f
C17 sky130_fd_pr__nfet_01v8_5Y6VJK_0.D vdd 0.0283f
C18 vin2 vin1 0.013356f
C19 vb2 Y 0.001182f
C20 vb2 vdd 0.028683f
C21 vb1 vin2 0.002591f
C22 sky130_fd_pr__nfet_01v8_5Y6VJK_0.D X 0.139332f
C23 vout2 vdd 8.10489f
C24 vb2 X 9.95e-19
C25 vout2 X 1.41382f
C26 sky130_fd_pr__nfet_01v8_DAKYLM_1.D vin1 3.04e-19
C27 vb2 sky130_fd_pr__nfet_01v8_5Y6VJK_0.D 0.062172f
C28 vout1 sky130_fd_pr__nfet_01v8_DAKYLM_1.D 0.773222f
C29 vb1 sky130_fd_pr__nfet_01v8_DAKYLM_1.D 0.174944f
C30 Y vin2 2.06e-19
C31 vin2 vdd 0.02161f
C32 sky130_fd_pr__nfet_01v8_5Y6VJK_0.D vout2 0.01051f
C33 vout1 vin1 1.34e-20
C34 vb1 vin1 0.006354f
C35 vb2 vout2 0.034526f
C36 vout1 vb1 0.001206f
C37 X vin2 0.033091f
C38 sky130_fd_pr__nfet_01v8_5Y6VJK_0.D vin2 0.014983f
C39 sky130_fd_pr__nfet_01v8_DAKYLM_1.D vdd 0.583158f
C40 sky130_fd_pr__nfet_01v8_DAKYLM_1.D Y 0.397725f
C41 vb2 vin2 0.001984f
C42 Y vin1 0.029862f
C43 vin1 vdd 0.020099f
C44 vout1 vdd 8.0091f
C45 vout1 Y 1.4029f
C46 X sky130_fd_pr__nfet_01v8_DAKYLM_1.D 4.16e-19
C47 vb1 Y 0.090448f
C48 vb1 vdd 0.323373f
C49 vout2 gnd 1.348106f
C50 vb2 gnd 0.977937f
C51 vin2 gnd 0.160939f
C52 vin1 gnd 0.161663f
C53 vb1 gnd 0.37867f
C54 vout1 gnd 2.024541f
C55 vdd gnd 18.239473f
C56 X gnd 1.663173f
C57 sky130_fd_pr__nfet_01v8_5Y6VJK_0.D gnd 0.554697f
C58 Y gnd 1.791587f
C59 sky130_fd_pr__nfet_01v8_DAKYLM_1.D gnd 7.0275f
C60 vout2.t8 gnd 0.519795f
C61 vout2.t5 gnd 0.143219f
C62 vout2.t2 gnd 0.143219f
C63 vout2.n0 gnd 0.313579f
C64 vout2.n1 gnd 1.44095f
C65 vout2.t10 gnd 0.143219f
C66 vout2.t6 gnd 0.143219f
C67 vout2.n2 gnd 0.313579f
C68 vout2.n3 gnd 0.697983f
C69 vout2.t3 gnd 0.143219f
C70 vout2.t1 gnd 0.143219f
C71 vout2.n4 gnd 0.313579f
C72 vout2.t7 gnd 0.143219f
C73 vout2.t4 gnd 0.143219f
C74 vout2.n5 gnd 0.313579f
C75 vout2.t0 gnd 0.103602f
C76 vout2.t9 gnd 0.489542f
C77 vout2.n6 gnd 0.594328f
C78 vout2.n7 gnd 0.797524f
C79 vout2.n8 gnd 0.697464f
C80 X.n0 gnd 0.209278f
C81 X.n1 gnd 0.233806f
C82 X.n2 gnd 0.23357f
C83 X.n3 gnd 0.072426f
C84 X.n4 gnd 0.167923f
C85 X.t8 gnd 0.095791f
C86 X.t11 gnd 0.095754f
C87 X.t6 gnd 0.095754f
C88 X.t10 gnd 0.095754f
C89 X.t4 gnd 0.095754f
C90 X.t7 gnd 0.095754f
C91 X.t2 gnd 0.095754f
C92 X.t9 gnd 0.095754f
C93 X.t5 gnd 0.095754f
C94 X.t3 gnd 0.095754f
C95 X.t1 gnd 0.031213f
C96 X.t0 gnd 0.085023f
C97 vdd.t1 gnd 0.069603f
C98 vdd.n0 gnd 0.044345f
C99 vdd.n1 gnd 0.065127f
C100 vdd.t38 gnd 1.19835f
C101 vdd.t32 gnd 0.437421f
C102 vdd.t26 gnd 0.437421f
C103 vdd.t42 gnd 0.437421f
C104 vdd.t34 gnd 0.328066f
C105 vdd.t39 gnd 0.054287f
C106 vdd.t33 gnd 0.054287f
C107 vdd.n2 gnd 0.159514f
C108 vdd.t31 gnd 0.054287f
C109 vdd.t41 gnd 0.054287f
C110 vdd.n3 gnd 0.161929f
C111 vdd.t25 gnd 0.054287f
C112 vdd.t37 gnd 0.054287f
C113 vdd.n4 gnd 0.159332f
C114 vdd.n5 gnd 0.396225f
C115 vdd.t35 gnd 0.054287f
C116 vdd.t29 gnd 0.054287f
C117 vdd.n6 gnd 0.159392f
C118 vdd.n7 gnd 0.198367f
C119 vdd.t27 gnd 0.054287f
C120 vdd.t43 gnd 0.054287f
C121 vdd.n8 gnd 0.159453f
C122 vdd.n9 gnd 0.204441f
C123 vdd.n10 gnd 0.27329f
C124 vdd.n11 gnd 0.47999f
C125 vdd.t28 gnd 0.328066f
C126 vdd.t24 gnd 0.437421f
C127 vdd.t36 gnd 0.437421f
C128 vdd.t30 gnd 0.437421f
C129 vdd.t40 gnd 1.09836f
C130 vdd.t0 gnd 0.915505f
C131 vdd.n12 gnd 0.392718f
C132 vdd.t23 gnd 0.069603f
C133 vdd.n13 gnd 0.044387f
C134 vdd.t12 gnd 1.19835f
C135 vdd.t8 gnd 0.437421f
C136 vdd.t16 gnd 0.437421f
C137 vdd.t20 gnd 0.437421f
C138 vdd.t6 gnd 0.328066f
C139 vdd.t2 gnd 1.19835f
C140 vdd.t10 gnd 0.437421f
C141 vdd.t4 gnd 0.437421f
C142 vdd.t18 gnd 0.437421f
C143 vdd.t14 gnd 0.328066f
C144 vdd.n14 gnd 0.47999f
C145 vdd.t13 gnd 0.054287f
C146 vdd.t9 gnd 0.054287f
C147 vdd.n15 gnd 0.161898f
C148 vdd.t11 gnd 0.054287f
C149 vdd.t3 gnd 0.054287f
C150 vdd.n16 gnd 0.162133f
C151 vdd.t19 gnd 0.054287f
C152 vdd.t5 gnd 0.054287f
C153 vdd.n17 gnd 0.159453f
C154 vdd.n18 gnd 0.400298f
C155 vdd.t7 gnd 0.054287f
C156 vdd.t15 gnd 0.054287f
C157 vdd.n19 gnd 0.159392f
C158 vdd.n20 gnd 0.198367f
C159 vdd.t17 gnd 0.054287f
C160 vdd.t21 gnd 0.054287f
C161 vdd.n21 gnd 0.159332f
C162 vdd.n22 gnd 0.190312f
C163 vdd.n23 gnd 0.243349f
C164 vdd.n24 gnd 0.090652f
C165 vdd.n25 gnd 0.093945f
C166 vdd.t22 gnd 0.815515f
C167 vdd.n26 gnd 0.392599f
C168 vout1.t0 gnd 0.134365f
C169 vout1.t9 gnd 0.134365f
C170 vout1.n0 gnd 0.294193f
C171 vout1.t6 gnd 0.134365f
C172 vout1.t4 gnd 0.134365f
C173 vout1.n1 gnd 0.294193f
C174 vout1.t10 gnd 0.097197f
C175 vout1.t2 gnd 0.459278f
C176 vout1.n2 gnd 0.593219f
C177 vout1.n3 gnd 0.74822f
C178 vout1.n4 gnd 0.654346f
C179 vout1.t5 gnd 0.48766f
C180 vout1.t3 gnd 0.134365f
C181 vout1.t7 gnd 0.134365f
C182 vout1.n5 gnd 0.294193f
C183 vout1.n6 gnd 1.35187f
C184 vout1.t8 gnd 0.134365f
C185 vout1.t1 gnd 0.134365f
C186 vout1.n7 gnd 0.294193f
C187 vout1.n8 gnd 0.654832f
C188 Y.n0 gnd 0.224762f
C189 Y.n1 gnd 0.251105f
C190 Y.n2 gnd 0.250851f
C191 Y.n3 gnd 0.077784f
C192 Y.n4 gnd 0.244018f
C193 Y.t6 gnd 0.102839f
C194 Y.t8 gnd 0.102878f
C195 Y.t2 gnd 0.102839f
C196 Y.t5 gnd 0.102839f
C197 Y.t10 gnd 0.102839f
C198 Y.t11 gnd 0.102839f
C199 Y.t7 gnd 0.102839f
C200 Y.t3 gnd 0.102839f
C201 Y.t9 gnd 0.102839f
C202 Y.t4 gnd 0.102839f
C203 Y.t0 gnd 0.033522f
C204 Y.t1 gnd 0.091314f
.ends

