magic
tech sky130A
magscale 1 2
timestamp 1720136304
<< error_p >>
rect -125 652 -67 658
rect 67 652 125 658
rect -125 618 -113 652
rect 67 618 79 652
rect -125 612 -67 618
rect 67 612 125 618
rect -221 -618 -163 -612
rect -29 -618 29 -612
rect 163 -618 221 -612
rect -221 -652 -209 -618
rect -29 -652 -17 -618
rect 163 -652 175 -618
rect -221 -658 -163 -652
rect -29 -658 29 -652
rect 163 -658 221 -652
<< pwell >>
rect -407 -790 407 790
<< nmos >>
rect -207 -580 -177 580
rect -111 -580 -81 580
rect -15 -580 15 580
rect 81 -580 111 580
rect 177 -580 207 580
<< ndiff >>
rect -269 568 -207 580
rect -269 -568 -257 568
rect -223 -568 -207 568
rect -269 -580 -207 -568
rect -177 568 -111 580
rect -177 -568 -161 568
rect -127 -568 -111 568
rect -177 -580 -111 -568
rect -81 568 -15 580
rect -81 -568 -65 568
rect -31 -568 -15 568
rect -81 -580 -15 -568
rect 15 568 81 580
rect 15 -568 31 568
rect 65 -568 81 568
rect 15 -580 81 -568
rect 111 568 177 580
rect 111 -568 127 568
rect 161 -568 177 568
rect 111 -580 177 -568
rect 207 568 269 580
rect 207 -568 223 568
rect 257 -568 269 568
rect 207 -580 269 -568
<< ndiffc >>
rect -257 -568 -223 568
rect -161 -568 -127 568
rect -65 -568 -31 568
rect 31 -568 65 568
rect 127 -568 161 568
rect 223 -568 257 568
<< psubdiff >>
rect -371 720 371 754
rect -371 -720 -337 720
rect 337 -720 371 720
rect -371 -754 -275 -720
rect 275 -754 371 -720
<< psubdiffcont >>
rect -275 -754 275 -720
<< poly >>
rect -129 652 -63 668
rect -129 618 -113 652
rect -79 618 -63 652
rect -207 580 -177 606
rect -129 602 -63 618
rect 63 652 129 668
rect 63 618 79 652
rect 113 618 129 652
rect -111 580 -81 602
rect -15 580 15 606
rect 63 602 129 618
rect 81 580 111 602
rect 177 580 207 606
rect -207 -602 -177 -580
rect -225 -618 -159 -602
rect -111 -606 -81 -580
rect -15 -602 15 -580
rect -225 -652 -209 -618
rect -175 -652 -159 -618
rect -225 -668 -159 -652
rect -33 -618 33 -602
rect 81 -606 111 -580
rect 177 -602 207 -580
rect -33 -652 -17 -618
rect 17 -652 33 -618
rect -33 -668 33 -652
rect 159 -618 225 -602
rect 159 -652 175 -618
rect 209 -652 225 -618
rect 159 -668 225 -652
<< polycont >>
rect -113 618 -79 652
rect 79 618 113 652
rect -209 -652 -175 -618
rect -17 -652 17 -618
rect 175 -652 209 -618
<< locali >>
rect -129 618 -113 652
rect -79 618 -63 652
rect 63 618 79 652
rect 113 618 129 652
rect -257 568 -223 584
rect -257 -584 -223 -568
rect -161 568 -127 584
rect -161 -584 -127 -568
rect -65 568 -31 584
rect -65 -584 -31 -568
rect 31 568 65 584
rect 31 -584 65 -568
rect 127 568 161 584
rect 127 -584 161 -568
rect 223 568 257 584
rect 223 -584 257 -568
rect -225 -652 -209 -618
rect -175 -652 -159 -618
rect -33 -652 -17 -618
rect 17 -652 33 -618
rect 159 -652 175 -618
rect 209 -652 225 -618
rect -291 -754 -275 -720
rect 275 -754 291 -720
<< viali >>
rect -113 618 -79 652
rect 79 618 113 652
rect -257 -568 -223 568
rect -161 -454 -127 454
rect -65 -568 -31 568
rect 31 -454 65 454
rect 127 -568 161 568
rect 223 -454 257 454
rect -209 -652 -175 -618
rect -17 -652 17 -618
rect 175 -652 209 -618
<< metal1 >>
rect -125 652 -67 658
rect -125 618 -113 652
rect -79 618 -67 652
rect -125 612 -67 618
rect 67 652 125 658
rect 67 618 79 652
rect 113 618 125 652
rect 67 612 125 618
rect -263 568 -217 580
rect -263 -568 -257 568
rect -223 -568 -217 568
rect -71 568 -25 580
rect -167 454 -121 466
rect -167 -454 -161 454
rect -127 -454 -121 454
rect -167 -466 -121 -454
rect -263 -580 -217 -568
rect -71 -568 -65 568
rect -31 -568 -25 568
rect 121 568 167 580
rect 25 454 71 466
rect 25 -454 31 454
rect 65 -454 71 454
rect 25 -466 71 -454
rect -71 -580 -25 -568
rect 121 -568 127 568
rect 161 -568 167 568
rect 217 454 263 466
rect 217 -454 223 454
rect 257 -454 263 454
rect 217 -466 263 -454
rect 121 -580 167 -568
rect -221 -618 -163 -612
rect -221 -652 -209 -618
rect -175 -652 -163 -618
rect -221 -658 -163 -652
rect -29 -618 29 -612
rect -29 -652 -17 -618
rect 17 -652 29 -618
rect -29 -658 29 -652
rect 163 -618 221 -612
rect 163 -652 175 -618
rect 209 -652 221 -618
rect 163 -658 221 -652
<< properties >>
string FIXED_BBOX -354 -737 354 737
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5.8 l 0.150 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 0 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 80 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
