magic
tech sky130A
magscale 1 2
timestamp 1756343927
<< error_p >>
rect -29 345 29 351
rect -29 311 -17 345
rect -29 305 29 311
<< nwell >>
rect -211 -484 211 484
<< pmos >>
rect -15 -336 15 264
<< pdiff >>
rect -73 252 -15 264
rect -73 -324 -61 252
rect -27 -324 -15 252
rect -73 -336 -15 -324
rect 15 252 73 264
rect 15 -324 27 252
rect 61 -324 73 252
rect 15 -336 73 -324
<< pdiffc >>
rect -61 -324 -27 252
rect 27 -324 61 252
<< nsubdiff >>
rect -175 414 175 448
rect -175 -414 -141 414
rect 141 -414 175 414
rect -175 -448 -79 -414
rect 79 -448 175 -414
<< nsubdiffcont >>
rect -79 -448 79 -414
<< poly >>
rect -33 345 33 361
rect -33 311 -17 345
rect 17 311 33 345
rect -33 295 33 311
rect -15 264 15 295
rect -15 -362 15 -336
<< polycont >>
rect -17 311 17 345
<< locali >>
rect -33 311 -17 345
rect 17 311 33 345
rect -61 252 -27 268
rect -61 -340 -27 -324
rect 27 252 61 268
rect 27 -340 61 -324
rect -95 -448 -79 -414
rect 79 -448 95 -414
<< viali >>
rect -17 311 17 345
rect -61 -324 -27 252
rect 27 -209 61 137
<< metal1 >>
rect -29 345 29 351
rect -29 311 -17 345
rect 17 311 29 345
rect -29 305 29 311
rect -67 252 -21 264
rect -67 -324 -61 252
rect -27 -324 -21 252
rect 21 137 67 149
rect 21 -209 27 137
rect 61 -209 67 137
rect 21 -221 67 -209
rect -67 -336 -21 -324
<< labels >>
rlabel nsubdiffcont 0 -431 0 -431 0 B
port 1 nsew
rlabel pdiffc -44 -36 -44 -36 0 D
port 2 nsew
rlabel pdiffc 44 -36 44 -36 0 S
port 3 nsew
rlabel polycont 0 328 0 328 0 G
port 4 nsew
<< properties >>
string FIXED_BBOX -158 -431 158 431
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 3 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 0 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 60 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1
<< end >>
