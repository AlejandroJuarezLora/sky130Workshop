magic
tech sky130A
magscale 1 2
timestamp 1734529318
<< pwell >>
rect -407 -790 407 790
<< nmos >>
rect -207 -580 -177 580
rect -111 -580 -81 580
rect -15 -580 15 580
rect 81 -580 111 580
rect 177 -580 207 580
<< ndiff >>
rect -269 568 -207 580
rect -269 -568 -257 568
rect -223 -568 -207 568
rect -269 -580 -207 -568
rect -177 568 -111 580
rect -177 -568 -161 568
rect -127 -568 -111 568
rect -177 -580 -111 -568
rect -81 568 -15 580
rect -81 -568 -65 568
rect -31 -568 -15 568
rect -81 -580 -15 -568
rect 15 568 81 580
rect 15 -568 31 568
rect 65 -568 81 568
rect 15 -580 81 -568
rect 111 568 177 580
rect 111 -568 127 568
rect 161 -568 177 568
rect 111 -580 177 -568
rect 207 568 269 580
rect 207 -568 223 568
rect 257 -568 269 568
rect 207 -580 269 -568
<< ndiffc >>
rect -257 -568 -223 568
rect -161 -568 -127 568
rect -65 -568 -31 568
rect 31 -568 65 568
rect 127 -568 161 568
rect 223 -568 257 568
<< psubdiff >>
rect -371 720 371 754
rect -371 -720 -337 720
rect 337 -720 371 720
rect -371 -754 -275 -720
rect 275 -754 371 -720
<< psubdiffcont >>
rect -275 -754 275 -720
<< poly >>
rect -129 652 -63 668
rect -129 618 -113 652
rect -79 618 -63 652
rect -207 580 -177 606
rect -129 602 -63 618
rect 63 652 129 668
rect 63 618 79 652
rect 113 618 129 652
rect -111 580 -81 602
rect -15 580 15 606
rect 63 602 129 618
rect 81 580 111 602
rect 177 580 207 606
rect -207 -602 -177 -580
rect -225 -618 -159 -602
rect -111 -606 -81 -580
rect -15 -602 15 -580
rect -225 -652 -209 -618
rect -175 -652 -159 -618
rect -225 -668 -159 -652
rect -33 -618 33 -602
rect 81 -606 111 -580
rect 177 -602 207 -580
rect -33 -652 -17 -618
rect 17 -652 33 -618
rect -33 -668 33 -652
rect 159 -618 225 -602
rect 159 -652 175 -618
rect 209 -652 225 -618
rect 159 -668 225 -652
<< polycont >>
rect -113 618 -79 652
rect 79 618 113 652
rect -209 -652 -175 -618
rect -17 -652 17 -618
rect 175 -652 209 -618
<< locali >>
rect -129 618 -113 652
rect -79 618 -63 652
rect 63 618 79 652
rect 113 618 129 652
rect -257 568 -223 584
rect -257 -584 -223 -568
rect -161 568 -127 584
rect -161 -584 -127 -568
rect -65 568 -31 584
rect -65 -584 -31 -568
rect 31 568 65 584
rect 31 -584 65 -568
rect 127 568 161 584
rect 127 -584 161 -568
rect 223 568 257 584
rect 223 -584 257 -568
rect -225 -652 -209 -618
rect -175 -652 -159 -618
rect -33 -652 -17 -618
rect 17 -652 33 -618
rect 159 -652 175 -618
rect 209 -652 225 -618
rect -291 -754 -275 -720
rect 275 -754 291 -720
<< viali >>
rect -113 618 -79 652
rect 79 618 113 652
rect -257 -568 -223 568
rect -161 -454 -127 454
rect -65 -568 -31 568
rect 31 -454 65 454
rect 127 -568 161 568
rect 223 -454 257 454
rect -209 -652 -175 -618
rect -17 -652 17 -618
rect 175 -652 209 -618
<< metal1 >>
rect -125 652 -67 658
rect 67 652 125 658
rect -125 618 -113 652
rect -79 618 79 652
rect 113 618 371 652
rect -125 612 -67 618
rect 67 612 125 618
rect -263 568 -217 580
rect -263 -568 -257 568
rect -223 -536 -217 568
rect -71 568 -25 580
rect -167 463 -121 466
rect -172 457 -120 463
rect -172 399 -161 405
rect -167 -454 -161 399
rect -127 399 -120 405
rect -127 -454 -121 399
rect -167 -466 -121 -454
rect -71 -536 -65 568
rect -223 -568 -65 -536
rect -31 -536 -25 568
rect 121 568 167 580
rect 25 464 71 466
rect 21 458 73 464
rect 21 400 31 406
rect 25 -454 31 400
rect 65 400 73 406
rect 65 -454 71 400
rect 25 -466 71 -454
rect 121 -536 127 568
rect -31 -568 127 -536
rect 161 -568 167 568
rect 217 465 263 466
rect 217 459 271 465
rect 217 407 219 459
rect 217 -454 223 407
rect 257 401 271 407
rect 257 -454 263 401
rect 217 -466 263 -454
rect -263 -569 167 -568
rect -263 -580 -217 -569
rect -71 -580 -25 -569
rect 121 -580 167 -569
rect -221 -618 -163 -612
rect -29 -618 29 -612
rect 163 -617 221 -612
rect 337 -617 371 618
rect 163 -618 371 -617
rect -221 -652 -209 -618
rect -175 -652 -17 -618
rect 17 -652 175 -618
rect 209 -651 371 -618
rect 209 -652 221 -651
rect -221 -658 -163 -652
rect -29 -658 29 -652
rect 163 -658 221 -652
<< via1 >>
rect -172 454 -120 457
rect -172 405 -161 454
rect -161 405 -127 454
rect -127 405 -120 454
rect 21 454 73 458
rect 21 406 31 454
rect 31 406 65 454
rect 65 406 73 454
rect 219 454 271 459
rect 219 407 223 454
rect 223 407 257 454
rect 257 407 271 454
<< metal2 >>
rect -178 448 -172 457
rect -327 413 -172 448
rect -178 405 -172 413
rect -120 449 -114 457
rect 15 449 21 458
rect -120 413 21 449
rect -120 405 -114 413
rect 15 406 21 413
rect 73 450 79 458
rect 213 450 219 459
rect 73 413 219 450
rect 73 406 79 413
rect 213 407 219 413
rect 271 407 277 459
<< labels >>
flabel metal1 s -101 -556 -101 -556 0 FreeSans 320 0 0 0 D
port 1 nsew
flabel metal2 s -327 413 -172 448 0 FreeSans 320 0 0 0 S
port 2 nsew
flabel locali s 8 -734 8 -734 0 FreeSans 320 0 0 0 B
port 3 nsew
flabel metal1 s 2 635 2 635 0 FreeSans 320 0 0 0 G
port 0 nsew
<< properties >>
string FIXED_BBOX -354 -737 354 737
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5.8 l 0.150 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 0 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 80 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
